module test2
  (
   /*AUTO-ARG*/
   INPUT             CLK,
   input wire        rst,
   
   input wire [31:0] in1,
   input WIRE        in2, in3,
   
   output wire       out1,
   output reg        out2, out3,
   
   inout             bidir1
   );



endmodule // test2
